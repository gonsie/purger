
module ccx ( cmp_gclk_c2_ccx_left, cmp_gclk_c2_ccx_right, scan_in, tcu_pce_ov, 
        gl_ccx_clk_stop_left, gl_ccx_clk_stop_right, tcu_aclk, tcu_bclk, 
        cpx_spc2_data_cx2, cpx_spc3_data_cx2, cpx_spc4_data_cx2, 
        cpx_spc5_data_cx2, cpx_spc6_data_cx2, cpx_spc7_data_cx2 );
  input [1:0] scan_in;
  output [1:0] scan_out;
  input [191:0] cpu_rep0_in;
  output [191:0] cpu_rep0_out;
  input [191:0] cpu_rep1_in;
  output [191:0] cpu_rep1_out;
  input [159:0] ccx_lstg_in;
  output [159:0] ccx_lstg_out;
  input [159:0] ccx_rstg_in;
  output [159:0] ccx_rstg_out;
  output [145:0] cpx_spc5_data_cx2;
  output [145:0] cpx_spc6_data_cx2;
  output [145:0] cpx_spc7_data_cx2;
  input cmp_gclk_c2_ccx_left, cmp_gclk_c2_ccx_right, tcu_pce_ov,
         gl_ccx_clk_stop_left, gl_ccx_clk_stop_right, tcu_aclk, tcu_bclk,
         tcu_scan_en, cluster_arst_l, tcu_atpg_mode, io_pcx_stall_pq,
         sctag0_pcx_stall_pq, sctag1_pcx_stall_pq, sctag2_pcx_stall_pq,
         sctag3_pcx_stall_pq, sctag4_pcx_stall_pq, sctag5_pcx_stall_pq,
         sctag6_pcx_stall_pq, sctag7_pcx_stall_pq, sctag0_cpx_atom_cq,
         sctag1_cpx_atom_cq, sctag2_cpx_atom_cq, sctag3_cpx_atom_cq,
         sctag4_cpx_atom_cq, sctag5_cpx_atom_cq, sctag6_cpx_atom_cq,
         sctag7_cpx_atom_cq;
  output pcx_fpio_data_rdy_px1, pcx_sctag0_atm_px1, pcx_sctag0_data_rdy_px1,
         pcx_sctag1_atm_px1, pcx_sctag1_data_rdy_px1, pcx_sctag2_atm_px1,
         pcx_sctag2_data_rdy_px1, pcx_sctag3_atm_px1, pcx_sctag3_data_rdy_px1,
         pcx_sctag4_atm_px1, pcx_sctag4_data_rdy_px1, pcx_sctag5_atm_px1,
         pcx_sctag5_data_rdy_px1, pcx_sctag6_atm_px1, pcx_sctag6_data_rdy_px1,
         pcx_sctag7_atm_px1, pcx_sctag7_data_rdy_px1;
  wire   \scan_in_buf[0] , tcu_pce_ov_buf, tcu_aclk_buf, tcu_bclk_buf,
         cluster_arst_l_buf, tcu_atpg_mode_buf, l2clk, tstgl_scan_out,
         clk_ccx_cclk_left, clk_ccx_cclk_right, cpx_sctag7_cpx_atom_rq_t,
         cpx_sctag6_cpx_atom_rq_t, cpx_sctag5_cpx_atom_rq_t,
         cpx_bfd2_i_dff_data_2_l1clk, cpx_bfd2_i_dff_data_3_l1clk,
         cpx_bfd3_i_dff_data_2_l1clk, cpx_bfd3_i_dff_data_3_l1clk,
         cpx_bfd4_i_dff_data_2_l1clk, cpx_bfd4_i_dff_data_3_l1clk,
         cpx_bfd5_i_dff_data_2_l1clk, cpx_bfd5_i_dff_data_3_l1clk,
         cpx_bfd6_i_dff_data_2_l1clk, cpx_bfd6_i_dff_data_3_l1clk,
         cpx_bfd7_i_dff_data_2_l1clk, cpx_bfd7_i_dff_data_3_l1clk,
         \pcx_arb8_qsel1_r_a[6] , \pcx_arb7_qsel1_r_a[6] ,
         \pcx_arb6_qsel1_r_a[6] , \pcx_arb5_qsel1_r_a[6] ,
         \pcx_arb4_qsel1_r_a[6] , \pcx_arb3_qsel1_r_a[6] ,
         \pcx_arb2_qsel1_r_a[6] , \pcx_arb1_qsel1_r_a[6] ,
         \pcx_arb0_qsel1_r_a[6] , pcx_sctag7_pcx_stall_pq_buf,
         pcx_sctag6_pcx_stall_pq_buf, pcx_sctag5_pcx_stall_pq_buf,
         pcx_sctag4_pcx_stall_pq_buf, pcx_sctag3_pcx_stall_pq_buf,
         pcx_pcx_arbl4_ard_stall_a_, pcx_pcx_arbl4_ard_fq_dir_a,
         n86382, n86383, n86384, n86385, n86386, n86387, n86388, n86389,
         n86390, n86391, n86392, n86393, n86394, n86395, n86396, n86397,
         n86398, n86399, n86400, n86401, n86402, n86403, n86404, n86405,
         n86406, n86407, n86408, n86409, n86410, n86411, n86412, n86413,
         n86414, n86415, n86416, n86417, n86418, n86419, n86420, n86421,
         n86422, n86423, n86424, n86425, n86426, n86427, n86428, n86429,
         n86430, n86431, n86432, n86433, n86434, n86435, n86436, n86437,
         n86438, n86439, n86440, n86441, n86442, n86443, n86444, n86445,
         n86446, n86447, n86448, n86449, n86450, n86451, n86452, n86453,
         n86454, n86455, n86456, n86457, n86458, n86459, n86460, n86461,
         n86462, n86463, n86464, n86465, n86466, n86467, n86468, n86469,
         n86470, n86471, n86472, n86473, n86474, n86475, n86476, n86477,
         n86478, n86479, n86480, n86481, n86482, n86483, n86484, n86485,
         n86486, n86487, n86488, n86489, n86490, n86491, n86492, n86493,
         n86494, n86495, n86496, n86497, n86498, n86499, n86500, n86501,
         n86502, n86503, n86504, n86505, n86506, n86507, n86508, n86509,
         n86510, n86511, n86512, n86513, n86514, n86515, n86516, n86517,
         n86518, n86519, n86520, n86521, n86522, n86523, n86524, n86525,
         n86526, n86527, n86528, n86529, n86530, n86531, n86532, n86533,
         n180675, n180676, n180677, n180678, n180679, n180680, n180681,
         n180682, n180683, n180684, n180685, n180686, n180687, n180688,
         n180689, n180690, n180691, n180692, n180693, n180694, n180695,
         n180696, n180697, n180698, n180699, n180700, n180701, n180702,
         n180703, n180704, n180705, n180706, n180707, n180708, n180709,
         n180710, n180711, n180712, n180713, n180714, n180715, n180716;
  wire   [7:0] cpx_io_cpx_req_rq;
  wire   [7:0] cpx_sctag7_cpx_req_rq;
  wire   [7:0] cpx_sctag6_cpx_req_rq;
  wire   [7:0] cpx_sctag5_cpx_req_rq;
  wire   [7:0] cpx_sctag4_cpx_req_rq;
  wire   [7:0] cpx_sctag3_cpx_req_rq;
  wire   [7:0] cpx_sctag2_cpx_req_rq;
  wire   [7:0] cpx_sctag1_cpx_req_rq;
  wire   [7:0] cpx_sctag0_cpx_req_rq;
  wire   [145:0] cpx_io_cpx_data_a_;
  wire   [7:0] cpx_io_cpx_req_cq_buf;
  wire   [145:0] cpx_io_cpx_data_ca_buf;
  wire   [7:5] cpx_cpx_dpa_cpx_dps0_arb_qsel1_r_a_rep;
  wire   [3:0] cpx_cpx_dpa_cpx_dps0_arb_qsel1_l_a_rep;
  wire   [4:2] cpx_cpx_arbr5_arc_add_281_carry;
  wire   [4:2] cpx_cpx_arbr5_arc_add_262_carry;
  wire   [4:2] cpx_cpx_arbr4_arc_add_281_carry;
  wire   [4:2] cpx_cpx_arbr4_arc_add_262_carry;
  wire   [4:2] cpx_cpx_arbl2_arc_add_262_carry;
  wire   [4:2] cpx_cpx_arbl1_arc_add_281_carry;
  wire   [4:2] cpx_cpx_arbl1_arc_add_262_carry;
  wire   [4:2] cpx_cpx_arbl0_arc_add_281_carry;
  wire   [4:2] cpx_cpx_arbl0_arc_add_262_carry;
  assign \scan_in_buf[0]  = scan_in[0];
  assign tcu_pce_ov_buf = tcu_pce_ov;
  assign tcu_aclk_buf = tcu_aclk;
  assign tcu_bclk_buf = tcu_bclk;
  assign cluster_arst_l_buf = cluster_arst_l;
  assign tcu_atpg_mode_buf = tcu_atpg_mode;
  assign cpx_sctag7_cpx_atom_rq_t = sctag7_cpx_atom_cq;
  assign cpx_sctag7_cpx_req_rq[7] = sctag7_cpx_req_cq[7];
  assign cpx_sctag7_cpx_req_rq[6] = sctag7_cpx_req_cq[6];
  assign cpx_sctag7_cpx_req_rq[5] = sctag7_cpx_req_cq[5];
  assign cpx_sctag7_cpx_req_rq[4] = sctag7_cpx_req_cq[4];
  assign cpx_sctag7_cpx_req_rq[3] = sctag7_cpx_req_cq[3];
  assign cpx_sctag7_cpx_req_rq[2] = sctag7_cpx_req_cq[2];
  assign cpx_sctag7_cpx_req_rq[1] = sctag7_cpx_req_cq[1];
  assign cpx_sctag7_cpx_req_rq[0] = sctag7_cpx_req_cq[0];
  assign cpx_sctag6_cpx_atom_rq_t = sctag6_cpx_atom_cq;
  assign cpx_sctag6_cpx_req_rq[7] = sctag6_cpx_req_cq[7];
  assign pcx_spc2_pcx_data_a[79] = spc2_pcx_data_pa[79];
  assign pcx_spc2_pcx_data_a[78] = spc2_pcx_data_pa[78];
  assign pcx_spc2_pcx_data_a[77] = spc2_pcx_data_pa[77];
  assign pcx_spc2_pcx_data_a[76] = spc2_pcx_data_pa[76];
  assign pcx_spc2_pcx_data_a[75] = spc2_pcx_data_pa[75];
  assign pcx_spc2_pcx_data_a[74] = spc2_pcx_data_pa[74];
  assign pcx_spc2_pcx_data_a[73] = spc2_pcx_data_pa[73];
  assign pcx_spc2_pcx_data_a[72] = spc2_pcx_data_pa[72];
  assign pcx_spc2_pcx_data_a[71] = spc2_pcx_data_pa[71];
  assign pcx_spc2_pcx_data_a[70] = spc2_pcx_data_pa[70];
  assign pcx_spc2_pcx_data_a[69] = spc2_pcx_data_pa[69];
  assign pcx_sctag6_pcx_stall_pq_buf = sctag6_pcx_stall_pq;
  assign pcx_sctag5_pcx_stall_pq_buf = sctag5_pcx_stall_pq;
  assign pcx_sctag4_pcx_stall_pq_buf = sctag4_pcx_stall_pq;
  assign pcx_sctag3_pcx_stall_pq_buf = sctag3_pcx_stall_pq;
  assign pcx_sctag2_pcx_stall_pq_buf = sctag2_pcx_stall_pq;
  assign pcx_sctag1_pcx_stall_pq_buf = sctag1_pcx_stall_pq;
  assign pcx_sctag0_pcx_stall_pq_buf = sctag0_pcx_stall_pq;
  assign pcx_io_pcx_stall_pq_buf = io_pcx_stall_pq;
  assign pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused = tcu_scan_en;
  assign pcx_spc5_grant_px[0] = pcx_pcx_dpa_pcx_dps0_pcx_rep_scan_rep3_out;

  n2_clk_ccx_cmp_cust clk_ccx_xtop ( .cclk_left(clk_ccx_cclk_left), 
        .cclk_right(clk_ccx_cclk_right), .l2clk(n138) );
  n2_clk_ccx_cmp_cust clk_ccx_xbottom ( .cclk_left(clk_ccx_cclk_left), 
        .cclk_right(clk_ccx_cclk_right), .l2clk(n139) );
  n2_clk_clstr_hdr_cust clk_ccx_xcluster_header_left ( .gclk(
        cmp_gclk_c2_ccx_left), .l2clk(l2clk), .cluster_arst_l(
        cluster_arst_l_buf), .ccu_div_ph(1'b1), .cluster_div_en(1'b0), 
        .tcu_div_bypass(1'b0), .scan_in(1'b0), .scan_en(1'b0), .tcu_aclk(1'b0), 
        .tcu_bclk(1'b0), .ccu_cmp_slow_sync_en(1'b0), .ccu_slow_cmp_sync_en(
        1'b0), .tcu_pce_ov(1'b1), .tcu_clk_stop(gl_ccx_clk_stop_left), 
        .rst_por_(1'b0), .rst_wmr_(1'b0), .rst_wmr_protect(1'b0), 
        .tcu_wr_inhibit(1'b0), .tcu_atpg_mode(tcu_atpg_mode_buf), .cclk(
        clk_ccx_cclk_left) );
  n2_clk_clstr_hdr_cust clk_ccx_xcluster_header_right ( .gclk(
        cmp_gclk_c2_ccx_right), .l2clk(l2clk), .cluster_arst_l(
        cluster_arst_l_buf), .ccu_div_ph(1'b1), .cluster_div_en(1'b0), 
        .tcu_div_bypass(1'b0), .scan_in(\scan_in_buf[0] ), .scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_aclk(tcu_aclk_buf), .tcu_bclk(tcu_bclk_buf), .ccu_cmp_slow_sync_en(1'b0), .ccu_slow_cmp_sync_en(
        1'b0), .tcu_pce_ov(tcu_pce_ov_buf), .tcu_clk_stop(
        gl_ccx_clk_stop_right), .rst_por_(1'b1), .rst_wmr_(1'b1), 
        .rst_wmr_protect(1'b0), .tcu_wr_inhibit(1'b0), .tcu_atpg_mode(
        tcu_atpg_mode_buf), .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), 
        .bclk(pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .cclk(
        clk_ccx_cclk_right) );
  n2_flop_bank_cust tstgl_i9 ( .l2clk(l2clk), .scan_in(tstgl_scan_out8), 
        .scan_out(tstgl_scan_out), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[159:144]), .data_in(ccx_lstg_in[159:144]) );
  n2_flop_bank_cust tstgl_i8 ( .l2clk(l2clk), .scan_in(tstgl_scan_out7), 
        .scan_out(tstgl_scan_out8), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[143:128]), .data_in(ccx_lstg_in[143:128]) );
  n2_flop_bank_cust tstgl_i7 ( .l2clk(l2clk), .scan_in(tstgl_scan_out6), 
        .scan_out(tstgl_scan_out7), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[127:112]), .data_in(ccx_lstg_in[127:112]) );
  n2_flop_bank_cust tstgl_i6 ( .l2clk(l2clk), .scan_in(tstgl_scan_out5), 
        .scan_out(tstgl_scan_out6), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[111:96]), .data_in(ccx_lstg_in[111:96]) );
  n2_flop_bank_cust tstgl_i5 ( .l2clk(l2clk), .scan_in(tstgl_scan_out4), 
        .scan_out(tstgl_scan_out5), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[95:80]), .data_in(ccx_lstg_in[95:80]) );
  n2_flop_bank_cust tstgl_i4 ( .l2clk(l2clk), .scan_in(tstgl_scan_out3), 
        .scan_out(tstgl_scan_out4), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[79:64]), .data_in(ccx_lstg_in[79:64]) );
  n2_flop_bank_cust tstgl_i3 ( .l2clk(l2clk), .scan_in(tstgl_scan_out2), 
        .scan_out(tstgl_scan_out3), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[63:48]), .data_in(ccx_lstg_in[63:48]) );
  n2_flop_bank_cust tstgl_i2 ( .l2clk(l2clk), .scan_in(tstgl_scan_out1), 
        .scan_out(tstgl_scan_out2), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[47:32]), .data_in(ccx_lstg_in[47:32]) );
  n2_flop_bank_cust tstgl_i1 ( .l2clk(l2clk), .scan_in(tstgl_scan_out0), 
        .scan_out(tstgl_scan_out1), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[31:16]), .data_in(ccx_lstg_in[31:16]) );
  n2_flop_bank_cust tstgl_i0 ( .l2clk(l2clk), .scan_in(
        pcx_pcx_dpa_pcx_dps6_pcx_mac7_i0_mac_c_q0[4]), .scan_out(
        tstgl_scan_out0), .tcu_aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_lstg_out[15:0]), .data_in(ccx_lstg_in[15:0]) );
  n2_flop_bank_cust tstgr_i9 ( .l2clk(l2clk), .scan_in(tstgr_scan_out8), 
        .scan_out(scan_out[1]), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[159:144]), .data_in(ccx_rstg_in[159:144]) );
  n2_flop_bank_cust tstgr_i8 ( .l2clk(l2clk), .scan_in(tstgr_scan_out7), 
        .scan_out(tstgr_scan_out8), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[143:128]), .data_in(ccx_rstg_in[143:128]) );
  n2_flop_bank_cust tstgr_i7 ( .l2clk(l2clk), .scan_in(tstgr_scan_out6), 
        .scan_out(tstgr_scan_out7), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[127:112]), .data_in(ccx_rstg_in[127:112]) );
  n2_flop_bank_cust tstgr_i6 ( .l2clk(l2clk), .scan_in(tstgr_scan_out5), 
        .scan_out(tstgr_scan_out6), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[111:96]), .data_in(ccx_rstg_in[111:96]) );
  n2_flop_bank_cust tstgr_i5 ( .l2clk(l2clk), .scan_in(tstgr_scan_out4), 
        .scan_out(tstgr_scan_out5), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[95:80]), .data_in(ccx_rstg_in[95:80]) );
  n2_flop_bank_cust tstgr_i4 ( .l2clk(l2clk), .scan_in(tstgr_scan_out3), 
        .scan_out(tstgr_scan_out4), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[79:64]), .data_in(ccx_rstg_in[79:64]) );
  n2_flop_bank_cust tstgr_i3 ( .l2clk(l2clk), .scan_in(tstgr_scan_out2), 
        .scan_out(tstgr_scan_out3), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[63:48]), .data_in(ccx_rstg_in[63:48]) );
  n2_flop_bank_cust tstgr_i2 ( .l2clk(l2clk), .scan_in(tstgr_scan_out1), 
        .scan_out(tstgr_scan_out2), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[47:32]), .data_in(ccx_rstg_in[47:32]) );
  n2_flop_bank_cust tstgr_i1 ( .l2clk(l2clk), .scan_in(tstgr_scan_out0), 
        .scan_out(tstgr_scan_out1), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[31:16]), .data_in(ccx_rstg_in[31:16]) );
  n2_flop_bank_cust tstgr_i0 ( .l2clk(l2clk), .scan_in(tstgl_scan_out), 
        .scan_out(tstgr_scan_out0), .tcu_aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .tcu_bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused), .tcu_scan_en(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .tcu_pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .local_stop(1'b0), 
        .data_out(ccx_rstg_out[15:0]), .data_in(ccx_rstg_in[15:0]) );
  AN4P U9592 ( .A(\pcx_pcx_arbr8_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr8_fifo_rptr_a[0]), .C(n83254), .D(n110199), .Z(n83253) );
  AN4P U9921 ( .A(\pcx_pcx_arbr7_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr7_fifo_rptr_a[0]), .C(n83548), .D(n110198), .Z(n83547) );
  AN4P U10250 ( .A(\pcx_pcx_arbr6_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr6_fifo_rptr_a[0]), .C(n83839), .D(n110197), .Z(n83838) );
  AN4P U10579 ( .A(\pcx_pcx_arbr5_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr5_fifo_rptr_a[0]), .C(n84130), .D(n110196), .Z(n84129) );
  AN4P U10908 ( .A(\pcx_pcx_arbr4_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr4_fifo_rptr_a[0]), .C(n84421), .D(n110195), .Z(n84420) );
  AN4P U11228 ( .A(\pcx_pcx_arbr3_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr3_fifo_rptr_a[0]), .C(n84697), .D(n110194), .Z(n84696) );
  AN4P U11548 ( .A(\pcx_pcx_arbr2_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr2_fifo_rptr_a[0]), .C(n84976), .D(n110193), .Z(n84975) );
  AN4P U11868 ( .A(\pcx_pcx_arbr1_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr1_fifo_rptr_a[0]), .C(n85255), .D(n110192), .Z(n85254) );
  AN4P U12188 ( .A(\pcx_pcx_arbr0_arc_rptr_a[4] ), .B(
        pcx_pcx_arbr0_fifo_rptr_a[0]), .C(n85534), .D(n110191), .Z(n85533) );
  AN4P U12508 ( .A(\pcx_pcx_arbl8_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl8_fifo_rptr_a[0]), .C(n85813), .D(n110190), .Z(n85812) );
  AN4P U12828 ( .A(\pcx_pcx_arbl7_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl7_fifo_rptr_a[0]), .C(n86092), .D(n110189), .Z(n86091) );
  AN4P U13148 ( .A(\pcx_pcx_arbl6_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl6_fifo_rptr_a[0]), .C(n86371), .D(n110188), .Z(n86370) );
  AN4P U13468 ( .A(\pcx_pcx_arbl5_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl5_fifo_rptr_a[0]), .C(n86650), .D(n110187), .Z(n86649) );
  AN4P U13788 ( .A(\pcx_pcx_arbl4_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl4_fifo_rptr_a[0]), .C(n86929), .D(n110186), .Z(n86928) );
  AN4P U14117 ( .A(\pcx_pcx_arbl3_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl3_fifo_rptr_a[0]), .C(n87223), .D(n110185), .Z(n87222) );
  AN4P U14446 ( .A(\pcx_pcx_arbl2_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl2_fifo_rptr_a[0]), .C(n87514), .D(n110184), .Z(n87513) );
  AN4P U14775 ( .A(\pcx_pcx_arbl1_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl1_fifo_rptr_a[0]), .C(n87805), .D(n110183), .Z(n87804) );
  AN4P U15104 ( .A(\pcx_pcx_arbl0_arc_rptr_a[4] ), .B(
        pcx_pcx_arbl0_fifo_rptr_a[0]), .C(n88096), .D(n110182), .Z(n88095) );
  AN4P U27517 ( .A(n88141), .B(n88131), .C(n97614), .D(n97615), .Z(n87902) );
  AN4P U27518 ( .A(n88150), .B(n88159), .C(n88168), .D(n88177), .Z(n97615) );
  AN4P U27852 ( .A(n83306), .B(n83317), .C(n83327), .D(n83338), .Z(n97751) );
  AO1P U28019 ( .A(n179229), .B(n108333), .C(n98051), .D(n98052), .Z(n98050)
         );
  AN2P U28098 ( .A(n98058), .B(n98088), .Z(n98093) );
  AN2P U28102 ( .A(pcx_pcx_arbl0_ard_stall_a_), .B(n169750), .Z(n98111) );
  AO1P U28115 ( .A(n179306), .B(n108331), .C(n98118), .D(n98119), .Z(n98117)
         );
  AN2P U28194 ( .A(n98125), .B(n98155), .Z(n98160) );
  AN2P U28198 ( .A(pcx_pcx_arbl1_ard_stall_a_), .B(n169638), .Z(n98178) );
  AO1P U28211 ( .A(n179383), .B(n108329), .C(n98185), .D(n98186), .Z(n98184)
         );
  AN2P U28290 ( .A(n98192), .B(n98222), .Z(n98227) );
  AN2P U28294 ( .A(pcx_pcx_arbl2_ard_stall_a_), .B(n169526), .Z(n98245) );
  AO1P U28307 ( .A(n179458), .B(n108327), .C(n98252), .D(n98253), .Z(n98251)
         );
  AN2P U28386 ( .A(n98259), .B(n98289), .Z(n98294) );
  AN2P U28390 ( .A(pcx_pcx_arbl3_ard_stall_a_), .B(n169414), .Z(n98312) );
  AO1P U29279 ( .A(n180217), .B(n180202), .C(n98861), .D(n98862), .Z(n98860)
         );
  AN2P U29358 ( .A(n98868), .B(n98898), .Z(n98903) );
  AN2P U29362 ( .A(pcx_pcx_arbr4_ard_stall_a_), .B(n168151), .Z(n98921) );
  AO1P U29375 ( .A(n180293), .B(n180278), .C(n98928), .D(n98929), .Z(n98927)
         );
  AN2P U29454 ( .A(n98935), .B(n98965), .Z(n98970) );
  AN2P U29458 ( .A(pcx_pcx_arbr5_ard_stall_a_), .B(n168039), .Z(n98988) );
  AO1P U29471 ( .A(n180369), .B(n180354), .C(n98995), .D(n98996), .Z(n98994)
         );
  AN2P U29550 ( .A(n99002), .B(n99032), .Z(n99037) );
  AN2P U29554 ( .A(pcx_pcx_arbr6_ard_stall_a_), .B(n167927), .Z(n99055) );
  AO1P U29567 ( .A(n180445), .B(n180430), .C(n99062), .D(n99063), .Z(n99061)
         );
  AN2P U29646 ( .A(n99069), .B(n99099), .Z(n99104) );
  AN2P U29650 ( .A(pcx_pcx_arbr7_ard_stall_a_), .B(n167815), .Z(n99122) );
  AN2P U29956 ( .A(n139), .B(n138), .Z(l2clk) );
  AN4P U40793 ( .A(\cpx_cpx_arbr7_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr7_fifo_rptr_a[0]), .C(n99599), .D(n110181), .Z(n99598) );
  AO1P U40948 ( .A(n108309), .B(n99422), .C(n99420), .D(n107319), .Z(
        cpx_cpx_arbr7_arc_input_req_sel_q) );
  AN2P U41022 ( .A(n99723), .B(n99725), .Z(n99716) );
  AN2P U41026 ( .A(cpx_cpx_arbr7_ard_stall_a_), .B(n169950), .Z(n99734) );
  AN4P U41038 ( .A(n99642), .B(n99632), .C(n99736), .D(n99737), .Z(n99421) );
  AN4P U41039 ( .A(n99653), .B(n99665), .C(n99677), .D(n99688), .Z(n99737) );
  AN4P U41252 ( .A(\cpx_cpx_arbr6_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr6_fifo_rptr_a[0]), .C(n99932), .D(n110180), .Z(n99931) );
  AO1P U41407 ( .A(n108307), .B(n99755), .C(n99753), .D(n107303), .Z(
        cpx_cpx_arbr6_arc_input_req_sel_q) );
  AN2P U41481 ( .A(n100056), .B(n100058), .Z(n100049) );
  AN2P U41485 ( .A(cpx_cpx_arbr6_ard_stall_a_), .B(n170097), .Z(n100067) );
  AN4P U41497 ( .A(n99975), .B(n99965), .C(n100069), .D(n100070), .Z(n99754)
         );
  AN4P U41498 ( .A(n99986), .B(n99998), .C(n100010), .D(n100021), .Z(n100070)
         );
  AN4P U41711 ( .A(\cpx_cpx_arbr5_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr5_fifo_rptr_a[0]), .C(n100265), .D(n110179), .Z(n100264)
         );
  AO1P U41866 ( .A(n108305), .B(n100088), .C(n100086), .D(n107287), .Z(
        cpx_cpx_arbr5_arc_input_req_sel_q) );
  AN2P U41940 ( .A(n100389), .B(n100391), .Z(n100382) );
  AN2P U41944 ( .A(cpx_cpx_arbr5_ard_stall_a_), .B(n170244), .Z(n100400) );
  AN4P U41956 ( .A(n100308), .B(n100298), .C(n100402), .D(n100403), .Z(n100087) );
  AN4P U41957 ( .A(n100319), .B(n100331), .C(n100343), .D(n100354), .Z(n100403) );
  AN4P U42170 ( .A(\cpx_cpx_arbr4_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr4_fifo_rptr_a[0]), .C(n100598), .D(n110178), .Z(n100597)
         );
  AO1P U42325 ( .A(n108303), .B(n100421), .C(n100419), .D(n107271), .Z(
        cpx_cpx_arbr4_arc_input_req_sel_q) );
  AN2P U42399 ( .A(n100722), .B(n100724), .Z(n100715) );
  AN2P U42403 ( .A(cpx_cpx_arbr4_ard_stall_a_), .B(n170391), .Z(n100733) );
  AN4P U42415 ( .A(n100641), .B(n100631), .C(n100735), .D(n100736), .Z(n100420) );
  AN4P U42416 ( .A(n100652), .B(n100664), .C(n100676), .D(n100687), .Z(n100736) );
  AN4P U42629 ( .A(\cpx_cpx_arbr3_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr3_fifo_rptr_a[0]), .C(n100931), .D(n110177), .Z(n100930)
         );
  AO1P U42784 ( .A(n108301), .B(n100754), .C(n100752), .D(n107255), .Z(
        cpx_cpx_arbr3_arc_input_req_sel_q) );
  AN2P U42858 ( .A(n101055), .B(n101057), .Z(n101048) );
  AN2P U42862 ( .A(cpx_cpx_arbr3_ard_stall_a_), .B(n170538), .Z(n101066) );
  AN4P U42874 ( .A(n100974), .B(n100964), .C(n101068), .D(n101069), .Z(n100753) );
  AN4P U42875 ( .A(n100985), .B(n100997), .C(n101009), .D(n101020), .Z(n101069) );
  AN4P U43088 ( .A(\cpx_cpx_arbr2_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr2_fifo_rptr_a[0]), .C(n101264), .D(n110176), .Z(n101263)
         );
  AO1P U43243 ( .A(n108299), .B(n101087), .C(n101085), .D(n107239), .Z(
        cpx_cpx_arbr2_arc_input_req_sel_q) );
  AN2P U43317 ( .A(n101388), .B(n101390), .Z(n101381) );
  AN2P U43321 ( .A(cpx_cpx_arbr2_ard_stall_a_), .B(n170687), .Z(n101399) );
  AN4P U43333 ( .A(n101307), .B(n101297), .C(n101401), .D(n101402), .Z(n101086) );
  AN4P U43334 ( .A(n101318), .B(n101330), .C(n101342), .D(n101353), .Z(n101402) );
  AN4P U43547 ( .A(\cpx_cpx_arbr1_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr1_fifo_rptr_a[0]), .C(n101597), .D(n110175), .Z(n101596)
         );
  AO1P U43702 ( .A(n108297), .B(n101420), .C(n101418), .D(n107223), .Z(
        cpx_cpx_arbr1_arc_input_req_sel_q) );
  AN2P U43776 ( .A(n101721), .B(n101723), .Z(n101714) );
  AN2P U43780 ( .A(cpx_cpx_arbr1_ard_stall_a_), .B(n170836), .Z(n101732) );
  AN4P U43792 ( .A(n101640), .B(n101630), .C(n101734), .D(n101735), .Z(n101419) );
  AN4P U43793 ( .A(n101651), .B(n101663), .C(n101675), .D(n101686), .Z(n101735) );
  AN4P U44006 ( .A(\cpx_cpx_arbr0_arc_rptr_a[4] ), .B(
        cpx_cpx_arbr0_fifo_rptr_a[0]), .C(n101930), .D(n110174), .Z(n101929)
         );
  AO1P U44161 ( .A(n108295), .B(n101753), .C(n101751), .D(n107207), .Z(
        cpx_cpx_arbr0_arc_input_req_sel_q) );
  AN2P U44235 ( .A(n102054), .B(n102056), .Z(n102047) );
  AN2P U44239 ( .A(cpx_cpx_arbr0_ard_stall_a_), .B(n170985), .Z(n102065) );
  AN4P U44251 ( .A(n101973), .B(n101963), .C(n102067), .D(n102068), .Z(n101752) );
  AN4P U44252 ( .A(n101984), .B(n101996), .C(n102008), .D(n102019), .Z(n102068) );
  AN4P U44465 ( .A(\cpx_cpx_arbl7_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl7_fifo_rptr_a[0]), .C(n102263), .D(n110173), .Z(n102262)
         );
  AO1P U44620 ( .A(n108293), .B(n102086), .C(n102084), .D(n107191), .Z(
        cpx_cpx_arbl7_arc_input_req_sel_q) );
  AN2P U44694 ( .A(n102385), .B(n102387), .Z(n102378) );
  AN2P U44698 ( .A(cpx_cpx_arbl7_ard_stall_a_), .B(n171092), .Z(n102396) );
  AN4P U44710 ( .A(n102312), .B(n102300), .C(n102398), .D(n102399), .Z(n102085) );
  AN4P U44711 ( .A(n102321), .B(n102331), .C(n102341), .D(n102350), .Z(n102399) );
  AN4P U44924 ( .A(\cpx_cpx_arbl6_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl6_fifo_rptr_a[0]), .C(n102594), .D(n110172), .Z(n102593)
         );
  AO1P U45079 ( .A(n108291), .B(n102417), .C(n102415), .D(n107175), .Z(
        cpx_cpx_arbl6_arc_input_req_sel_q) );
  AN2P U45153 ( .A(n102716), .B(n102718), .Z(n102709) );
  AN2P U45157 ( .A(cpx_cpx_arbl6_ard_stall_a_), .B(n171171), .Z(n102727) );
  AN4P U45169 ( .A(n102643), .B(n102631), .C(n102729), .D(n102730), .Z(n102416) );
  AN4P U45170 ( .A(n102652), .B(n102662), .C(n102672), .D(n102681), .Z(n102730) );
  AN4P U45383 ( .A(\cpx_cpx_arbl5_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl5_fifo_rptr_a[0]), .C(n102925), .D(n110171), .Z(n102924)
         );
  AO1P U45538 ( .A(n108289), .B(n102748), .C(n102746), .D(n107159), .Z(
        cpx_cpx_arbl5_arc_input_req_sel_q) );
  AN2P U45612 ( .A(n103047), .B(n103049), .Z(n103040) );
  AN2P U45616 ( .A(cpx_cpx_arbl5_ard_stall_a_), .B(n171250), .Z(n103058) );
  AN4P U45628 ( .A(n102974), .B(n102962), .C(n103060), .D(n103061), .Z(n102747) );
  AN4P U45629 ( .A(n102983), .B(n102993), .C(n103003), .D(n103012), .Z(n103061) );
  AN4P U45842 ( .A(\cpx_cpx_arbl4_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl4_fifo_rptr_a[0]), .C(n103256), .D(n110170), .Z(n103255)
         );
  AO1P U45997 ( .A(n108287), .B(n103079), .C(n103077), .D(n107143), .Z(
        cpx_cpx_arbl4_arc_input_req_sel_q) );
  AN2P U46071 ( .A(n103378), .B(n103380), .Z(n103371) );
  AN2P U46075 ( .A(cpx_cpx_arbl4_ard_stall_a_), .B(n171329), .Z(n103389) );
  AN4P U46087 ( .A(n103305), .B(n103293), .C(n103391), .D(n103392), .Z(n103078) );
  AN4P U46088 ( .A(n103314), .B(n103324), .C(n103334), .D(n103343), .Z(n103392) );
  AN4P U46301 ( .A(\cpx_cpx_arbl3_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl3_fifo_rptr_a[0]), .C(n103587), .D(n110169), .Z(n103586)
         );
  AO1P U46456 ( .A(n108285), .B(n103410), .C(n103408), .D(n107127), .Z(
        cpx_cpx_arbl3_arc_input_req_sel_q) );
  AN2P U46530 ( .A(n103709), .B(n103711), .Z(n103702) );
  AN2P U46534 ( .A(cpx_cpx_arbl3_ard_stall_a_), .B(n171408), .Z(n103720) );
  AN4P U46546 ( .A(n103636), .B(n103624), .C(n103722), .D(n103723), .Z(n103409) );
  AN4P U46547 ( .A(n103645), .B(n103655), .C(n103665), .D(n103674), .Z(n103723) );
  AN4P U46760 ( .A(\cpx_cpx_arbl2_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl2_fifo_rptr_a[0]), .C(n103918), .D(n110168), .Z(n103917)
         );
  AO1P U46915 ( .A(n108283), .B(n103741), .C(n103739), .D(n107111), .Z(
        cpx_cpx_arbl2_arc_input_req_sel_q) );
  AN2P U46989 ( .A(n104040), .B(n104042), .Z(n104033) );
  AN2P U46993 ( .A(cpx_cpx_arbl2_ard_stall_a_), .B(n171487), .Z(n104051) );
  AN4P U47005 ( .A(n103967), .B(n103955), .C(n104053), .D(n104054), .Z(n103740) );
  AN4P U47006 ( .A(n103976), .B(n103986), .C(n103996), .D(n104005), .Z(n104054) );
  AN4P U47219 ( .A(\cpx_cpx_arbl1_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl1_fifo_rptr_a[0]), .C(n104249), .D(n110167), .Z(n104248)
         );
  AO1P U47374 ( .A(n108281), .B(n104072), .C(n104070), .D(n107095), .Z(
        cpx_cpx_arbl1_arc_input_req_sel_q) );
  AN2P U47448 ( .A(n104371), .B(n104373), .Z(n104364) );
  AN2P U47452 ( .A(cpx_cpx_arbl1_ard_stall_a_), .B(n171566), .Z(n104382) );
  AN4P U47464 ( .A(n104298), .B(n104286), .C(n104384), .D(n104385), .Z(n104071) );
  AN4P U47465 ( .A(n104307), .B(n104317), .C(n104327), .D(n104336), .Z(n104385) );
  AN4P U47678 ( .A(\cpx_cpx_arbl0_arc_rptr_a[4] ), .B(
        cpx_cpx_arbl0_fifo_rptr_a[0]), .C(n104580), .D(n110166), .Z(n104579)
         );
  AO1P U47833 ( .A(n108279), .B(n104403), .C(n104401), .D(n107079), .Z(
        cpx_cpx_arbl0_arc_input_req_sel_q) );
  AN2P U47907 ( .A(n104702), .B(n104704), .Z(n104695) );
  AN2P U47911 ( .A(cpx_cpx_arbl0_ard_stall_a_), .B(n171645), .Z(n104713) );
  AN4P U47923 ( .A(n104629), .B(n104617), .C(n104715), .D(n104716), .Z(n104402) );
  AN4P U47924 ( .A(n104638), .B(n104648), .C(n104658), .D(n104667), .Z(n104716) );
  OR3 U75332 ( .A(n167703), .B(n107544), .C(n83075), .Z(n83074) );
  OR3 U75333 ( .A(n167703), .B(n83075), .C(n83246), .Z(n83240) );
  OR3 U75334 ( .A(n167815), .B(n107537), .C(n83354), .Z(n83353) );
  OR3 U75335 ( .A(n83356), .B(n83357), .C(n83358), .Z(
        pcx_pcx_arbr7_ard_i_nor_atom_d0_0_N1) );
  OR3 U75336 ( .A(n167815), .B(n83354), .C(n83540), .Z(n83534) );
  OR3 U75337 ( .A(n167927), .B(n107529), .C(n83645), .Z(n83644) );
  OR3 U75338 ( .A(n83647), .B(n83648), .C(n83649), .Z(
        pcx_pcx_arbr6_ard_i_nor_atom_d0_0_N1) );
  OR3 U75339 ( .A(n167927), .B(n83645), .C(n83831), .Z(n83825) );
  OR3 U75340 ( .A(n168039), .B(n107521), .C(n83936), .Z(n83935) );
  OR3 U75341 ( .A(n83938), .B(n83939), .C(n83940), .Z(
        pcx_pcx_arbr5_ard_i_nor_atom_d0_0_N1) );
  OR3 U75342 ( .A(n168039), .B(n83936), .C(n84122), .Z(n84116) );
  OR3 U75343 ( .A(n168151), .B(n107513), .C(n84227), .Z(n84226) );
  OR3 U75344 ( .A(n84229), .B(n84230), .C(n84231), .Z(
        pcx_pcx_arbr4_ard_i_nor_atom_d0_0_N1) );
  OR3 U75345 ( .A(n168151), .B(n84227), .C(n84413), .Z(n84407) );
  OR3 U75363 ( .A(n169341), .B(n86750), .C(n86921), .Z(n86915) );
  OR3 U75364 ( .A(n169414), .B(n107360), .C(n87029), .Z(n87028) );
  OR3 U75365 ( .A(n87031), .B(n87032), .C(n87033), .Z(
        pcx_pcx_arbl3_ard_i_nor_atom_d0_0_N1) );
  OR3 U75366 ( .A(n169414), .B(n87029), .C(n87215), .Z(n87209) );
  OR3 U75367 ( .A(n169526), .B(n107352), .C(n87320), .Z(n87319) );
  OR3 U75368 ( .A(n87322), .B(n87323), .C(n87324), .Z(
        pcx_pcx_arbl2_ard_i_nor_atom_d0_0_N1) );
  OR3 U75369 ( .A(n169526), .B(n87320), .C(n87506), .Z(n87500) );
  OR3 U75370 ( .A(n169638), .B(n107344), .C(n87611), .Z(n87610) );
  OR3 U75371 ( .A(n87613), .B(n87614), .C(n87615), .Z(
        pcx_pcx_arbl1_ard_i_nor_atom_d0_0_N1) );
  OR3 U75372 ( .A(n169638), .B(n87611), .C(n87797), .Z(n87791) );
  OR3 U75373 ( .A(n169750), .B(n107336), .C(n87902), .Z(n87901) );
  OR3 U75374 ( .A(n87904), .B(n87905), .C(n87906), .Z(
        pcx_pcx_arbl0_ard_i_nor_atom_d0_0_N1) );
  OR3 U75375 ( .A(n169750), .B(n87902), .C(n88088), .Z(n88082) );
  OR3 U75399 ( .A(n83499), .B(n83481), .C(n83516), .Z(n83356) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[0]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[0]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[0]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[1]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[1]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[1]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[2]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[2]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[2]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[3]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[3]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[3]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[4]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[4]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[4]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[5]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[5]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[5]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[6]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[6]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[6]) );
  FD1 \cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_msff0_q_reg[7]  ( .D(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0_in[7]), .CP(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_l1clk0), .Q(
        cpx_cpx_dpa_cpx_dps0_cpx_mac0_i0_mac_b_q0[7]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem2_d0_0_q_reg[7]  ( .D(n178051), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata2[7]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem1_d0_0_q_reg[7]  ( .D(n178051), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata1[7]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem0_d0_0_q_reg[7]  ( .D(n178051), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata0[7]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_reqreg_d0_0_q_reg[7]  ( .D(
        cpx_cpx_arbl0_ard_fq_req[7]), .CP(cpx_cpx_arbl0_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl0_ard_fq_req_a[7]) );
  FD1 \cpx_cpx_arbl0_arc_q8_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178053), .CP(
        cpx_cpx_arbl0_arc_l1clk), .Q(cpx_cpx_arbl0_qfullbar_a[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem17_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata17[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem16_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata16[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem15_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata15[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem14_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata14[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem13_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata13[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem12_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata12[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem11_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata11[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem10_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata10[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem9_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata9[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem8_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata8[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem7_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata7[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem6_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata6[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem5_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata5[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem4_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata4[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem3_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata3[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem2_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata2[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem1_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata1[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem0_d0_0_q_reg[8]  ( .D(n178055), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata0[8]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_reqreg_d0_0_q_reg[8]  ( .D(
        cpx_cpx_arbl0_ard_fq_req[8]), .CP(cpx_cpx_arbl0_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl0_ard_fq_req_a[8]) );
  FD1 \cpx_cpx_arbl0_arc_q0_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178021), .CP(
        cpx_cpx_arbl0_arc_l1clk), .Q(cpx_cpx_arbl0_qfullbar_a[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem17_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata17[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem16_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata16[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem15_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata15[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem14_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata14[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem13_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata13[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem12_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata12[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem11_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata11[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem10_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata10[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem9_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata9[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem8_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata8[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem7_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata7[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem6_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata6[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem5_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata5[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem4_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata4[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem3_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata3[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem2_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata2[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem1_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata1[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_fmem0_d0_0_q_reg[0]  ( .D(n178023), .CP(
        cpx_cpx_arbl0_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl0_ard_fifo_rdata0[0]) );
  FD1 \cpx_cpx_arbl0_ard_i_dff_reqreg_d0_0_q_reg[0]  ( .D(
        cpx_cpx_arbl0_ard_fq_req[0]), .CP(cpx_cpx_arbl0_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl0_ard_fq_req_a[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_atom_a_d0_0_q_reg[9]  ( .D(n130396), .CP(
        cpx_cpx_arbl1_ard_i_dff_atom_a_l1clk), .Q(cpx_cpx_arbl1_ard_dir_a_) );
  FD1 \cpx_cpx_arbl1_arc_q4_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178111), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[4]) );
  FD1 \cpx_cpx_arbl1_arc_q3_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178107), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[3]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[3]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[3]) );
  FD1 \cpx_cpx_arbl1_arc_q1_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178099), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[1]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[1]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[9]  ( .D(n171568), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[9]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[1]  ( .D(n178101), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[1]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[2]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[2]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[2]) );
  FD1 \cpx_cpx_arbl1_arc_q2_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178103), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[2]  ( .D(n178105), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[2]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[3]  ( .D(n178109), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[3]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[4]  ( .D(n178113), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[4]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[4]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[4]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[9]  ( .D(n171569), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[9]) );
  FD1 \cpx_cpx_arbl1_arc_q5_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178115), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[5]  ( .D(n178117), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[5]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[5]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[5]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[5]) );
  FD1 \cpx_cpx_arbl1_arc_q6_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178119), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[6]  ( .D(n178121), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[6]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[6]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[6]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[6]) );
  FD1 \cpx_cpx_arbl1_arc_q7_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178123), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[7]  ( .D(n178125), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[7]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[7]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[7]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[7]) );
  FD1 \cpx_cpx_arbl1_arc_q8_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178127), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[8]  ( .D(n178129), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[8]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[8]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[8]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[8]) );
  FD1 \cpx_cpx_arbl1_arc_q0_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178095), .CP(
        cpx_cpx_arbl1_arc_l1clk), .Q(cpx_cpx_arbl1_qfullbar_a[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem17_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata17[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem16_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem16_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata16[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem15_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem15_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata15[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem14_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata14[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem13_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata13[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem12_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem12_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata12[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem11_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem11_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata11[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem10_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata10[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem9_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata9[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem8_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata8[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem7_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem7_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata7[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem6_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata6[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem5_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata5[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem4_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata4[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem3_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem3_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata3[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem2_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata2[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem1_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem1_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata1[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_fmem0_d0_0_q_reg[0]  ( .D(n178097), .CP(
        cpx_cpx_arbl1_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl1_ard_fifo_rdata0[0]) );
  FD1 \cpx_cpx_arbl1_ard_i_dff_reqreg_d0_0_q_reg[0]  ( .D(
        cpx_cpx_arbl1_ard_fq_req[0]), .CP(cpx_cpx_arbl1_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl1_ard_fq_req_a[0]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_atom_a_d0_0_q_reg[9]  ( .D(n130395), .CP(
        cpx_cpx_arbl2_ard_i_dff_atom_a_l1clk), .Q(cpx_cpx_arbl2_ard_dir_a_) );
  FD1 \cpx_cpx_arbl2_arc_q4_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178185), .CP(
        cpx_cpx_arbl2_arc_l1clk), .Q(cpx_cpx_arbl2_qfullbar_a[4]) );
  FD1 \cpx_cpx_arbl2_arc_q3_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178181), .CP(
        cpx_cpx_arbl2_arc_l1clk), .Q(cpx_cpx_arbl2_qfullbar_a[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_reqreg_d0_0_q_reg[3]  ( .D(
        cpx_cpx_arbl2_ard_fq_req[3]), .CP(cpx_cpx_arbl2_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl2_ard_fq_req_a[3]) );
  FD1 \cpx_cpx_arbl2_arc_q1_dff_qfullbar_a_d0_0_q_reg[0]  ( .D(n178173), .CP(
        cpx_cpx_arbl2_arc_l1clk), .Q(cpx_cpx_arbl2_qfullbar_a[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_reqreg_d0_0_q_reg[1]  ( .D(
        cpx_cpx_arbl2_ard_fq_req[1]), .CP(cpx_cpx_arbl2_ard_i_dff_reqreg_l1clk), .Q(cpx_cpx_arbl2_ard_fq_req_a[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem9_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata9[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem9_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata9[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem9_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata9[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem9_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem9_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata9[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem4_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata4[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem4_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata4[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem4_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata4[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem4_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem4_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata4[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem13_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata13[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem13_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata13[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem13_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata13[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem13_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem13_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata13[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem6_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata6[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem6_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata6[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem6_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata6[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem6_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem6_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata6[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem2_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata2[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem2_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata2[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem2_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata2[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem2_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem2_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata2[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem14_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata14[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem14_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata14[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem14_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata14[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem14_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem14_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata14[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem10_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata10[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem10_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata10[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem10_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata10[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem10_d0_0_q_reg[9]  ( .D(n171489), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem10_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata10[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem0_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata0[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem0_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata0[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem0_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata0[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem0_d0_0_q_reg[9]  ( .D(n171490), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem0_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata0[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem17_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata17[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem17_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata17[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem17_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata17[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem17_d0_0_q_reg[9]  ( .D(n171490), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem17_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata17[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem8_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata8[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem8_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata8[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem8_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata8[4]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem8_d0_0_q_reg[9]  ( .D(n171490), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem8_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata8[9]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem5_d0_0_q_reg[1]  ( .D(n178175), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata5[1]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem5_d0_0_q_reg[3]  ( .D(n178183), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata5[3]) );
  FD1 \cpx_cpx_arbl2_ard_i_dff_fmem5_d0_0_q_reg[4]  ( .D(n178187), .CP(
        cpx_cpx_arbl2_ard_i_dff_fmem5_l1clk), .Q(
        cpx_cpx_arbl2_ard_fifo_rdata5[4]) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps7_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107760), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps7_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107760), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps7_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107760), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps7_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac6_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac6_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107760), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb7_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps7_pcx_mac7_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps7_pcx_mac7_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107764), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac0_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac0_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107696), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac1_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac1_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107700), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac2_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac2_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107698), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_l_a_rep[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac3_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac3_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107702), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[5]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac4_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac4_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107770), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep_7), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac5_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac5_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107774), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_dpa_pcx_dps8_arb_qsel1_r_a_rep[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac6_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac6_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107768), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i0_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i0_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i0_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i0_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i1_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i1_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i1_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i1_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i2_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i2_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i2_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i2_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i3_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i3_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i3_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i3_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i4_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i4_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i4_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i4_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i5_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i5_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i5_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i5_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i6_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i6_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i6_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i6_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i7_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i7_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i7_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i7_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i8_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i8_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i8_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i8_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i9_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i9_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i9_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i9_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i10_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i10_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i10_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i10_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i11_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i11_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i11_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i11_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i12_c0_hdr1 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i12_l1clk1), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        \pcx_arb8_qsel1_r_a[6] ), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_ccx_l1hdr_16x pcx_pcx_dpa_pcx_dps8_pcx_mac7_i12_c0_hdr0 ( .l1clk(
        pcx_pcx_dpa_pcx_dps8_pcx_mac7_i12_l1clk0), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(n107772), 
        .pce_ov(pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), 
        .aclk(pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd_io_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd_io_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd0_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd0_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd1_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd1_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd2_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd2_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd3_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd3_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd4_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd4_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd5_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd5_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd6_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd6_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd7_i_dff_data_0_c0_0 ( .l1clk(
        pcx_bfd7_i_dff_data_0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd_io_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd_io_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd0_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd0_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd1_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd1_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd2_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd2_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd3_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd3_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd4_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd4_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd5_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd5_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd6_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd6_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd7_i_dff_data_1_c0_0 ( .l1clk(
        pcx_bfd7_i_dff_data_1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd_io_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd_io_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd_io_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd_io_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd0_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd0_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd0_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd0_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd1_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd1_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd1_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd1_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd2_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd2_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd2_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd2_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd3_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd3_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd3_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd3_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd4_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd4_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd4_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd4_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd5_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd5_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd5_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd5_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd6_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd6_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd6_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd6_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd7_i_dff_data_2_c0_0 ( .l1clk(
        pcx_bfd7_i_dff_data_2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_bfd7_i_dff_data_3_c0_0 ( .l1clk(
        pcx_bfd7_i_dff_data_3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl0_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl0_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl1_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl1_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl2_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl2_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl3_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl3_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl4_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl4_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl5_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl5_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl6_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl6_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbl7_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbl7_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr0_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr0_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr1_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr1_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr2_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr2_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr3_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr3_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr4_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr4_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr5_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr5_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr6_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr6_arc_l1clk) );
  cl_sc1_l1hdr_8x cpx_cpx_arbr7_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        cpx_cpx_arbr7_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl0_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl0_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl1_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl1_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl2_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl2_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl3_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl3_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl4_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl4_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl5_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl5_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl6_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl6_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl7_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl7_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbl8_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbl8_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr0_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr0_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr1_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr1_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr2_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr2_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr3_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr3_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr4_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr4_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr5_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr5_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr6_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr6_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr7_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr7_arc_l1clk) );
  cl_sc1_l1hdr_8x pcx_pcx_arbr8_arc_clkgen_c_0 ( .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .l1clk(
        pcx_pcx_arbr8_arc_l1clk) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl1_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl1_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl1_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl1_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl2_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl2_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl2_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl2_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl3_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl3_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl3_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl3_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl4_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl4_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl4_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl4_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl5_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl5_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl5_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl5_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl6_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl6_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl6_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl6_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl7_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbl7_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl7_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbl7_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr0_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr0_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr0_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr0_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr1_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr1_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr1_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr1_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr2_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr2_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr2_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr2_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr3_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr3_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr3_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr3_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr4_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr4_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr4_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr4_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr5_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr5_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr5_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr5_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr6_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr6_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr6_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr6_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr7_ard_i_dff_atom_a_c0_0 ( .l1clk(
        cpx_cpx_arbr7_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbr7_ard_i_dff_req_a_c0_0 ( .l1clk(
        cpx_cpx_arbr7_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl0_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl0_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl0_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl0_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl1_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl1_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl1_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl1_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl2_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl2_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl2_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl2_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl3_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl3_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl3_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl3_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl4_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl4_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl4_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl4_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl5_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl5_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl5_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl5_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl6_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl6_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl6_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl6_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl7_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl7_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl7_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl7_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl8_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbl8_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbl8_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbl8_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr0_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr0_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr0_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr0_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr1_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr1_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr1_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr1_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr2_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr2_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr2_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr2_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr3_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr3_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr3_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr3_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr4_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr4_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr4_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr4_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr5_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr5_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr5_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr5_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr6_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr6_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr6_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr6_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr7_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr7_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr7_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr7_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_atom_a_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_atom_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_req_a_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_req_a_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_penc2_8x cpx_cpx_arbl0_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl0_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl0_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl0_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl1_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl1_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl1_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl1_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl2_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl2_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl2_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl2_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl3_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl3_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl3_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl3_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl4_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl4_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl4_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl4_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl5_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl5_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl5_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl5_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl6_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl6_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl6_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl6_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl7_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbl7_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbl7_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbl7_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr0_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr0_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr0_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr0_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr1_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr1_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr1_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr1_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr2_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr2_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr2_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr2_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr3_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr3_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr3_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr3_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr4_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr4_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr4_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr4_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr5_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr5_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr5_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr5_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr6_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr6_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr6_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr6_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbr7_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        cpx_cpx_arbr7_fifo_rptr_a[0]), .psel0(
        cpx_cpx_arbr7_ard_i_mux_fmem17_16_psel0), .psel1(
        cpx_cpx_arbr7_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl0_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl0_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl0_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl0_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl1_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl1_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl1_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl1_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl2_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl2_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl2_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl2_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl3_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl3_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl3_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl3_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl4_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl4_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl4_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl4_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl5_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl5_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl5_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl5_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl6_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl6_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl6_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl6_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl7_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl7_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl7_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl7_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbl8_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbl8_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbl8_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbl8_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr0_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr0_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr0_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr0_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr1_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr1_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr1_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr1_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr2_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr2_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr2_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr2_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr3_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr3_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr3_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr3_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr4_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr4_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr4_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr4_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr5_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr5_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr5_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr5_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr6_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr6_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr6_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr6_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr7_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr7_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr7_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr7_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr8_ard_i_mux_fmem17_16_c0_0 ( .sel0(
        pcx_pcx_arbr8_fifo_rptr_a[0]), .psel0(
        pcx_pcx_arbr8_ard_i_mux_fmem17_16_psel0), .psel1(
        pcx_pcx_arbr8_ard_i_mux_fmem17_16_psel1) );
  cl_dp1_pdec8_8x cpx_cpx_arbl0_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl0_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl0_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl0_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl0_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl0_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl0_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl0_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl1_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl1_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl1_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl1_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl1_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl1_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl1_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl1_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl2_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl2_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl2_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl2_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl2_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl2_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl2_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl2_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl3_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl3_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl3_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl3_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl3_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl3_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl3_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl3_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl4_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl4_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl4_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl4_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl4_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl4_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl4_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl4_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl5_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl5_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl5_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl5_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl5_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl5_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl5_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl5_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl6_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl6_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl6_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl6_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl6_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl6_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl6_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl6_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl7_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbl7_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl7_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbl7_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbl7_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbl7_fifo_rptr_a[0]), .sel1(cpx_cpx_arbl7_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbl7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbl7_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr0_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr0_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr0_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr0_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr0_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr0_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr0_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr0_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr1_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr1_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr1_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr1_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr1_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr1_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr1_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr1_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr2_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr2_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr2_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr2_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr2_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr2_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr2_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr2_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr3_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr3_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr3_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr3_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr3_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr3_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr3_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr3_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr4_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr4_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr4_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr4_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr4_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr4_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr4_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr4_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr5_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr5_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr5_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr5_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr5_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr5_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr5_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr5_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr6_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr6_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr6_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr6_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr6_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr6_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr6_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr6_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr7_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        cpx_cpx_arbr7_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr7_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel0), .psel1(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel1), .psel2(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel2), .psel3(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel3), .psel4(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel4), .psel5(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel5), .psel6(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel6), .psel7(
        cpx_cpx_arbr7_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x cpx_cpx_arbr7_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        cpx_cpx_arbr7_fifo_rptr_a[0]), .sel1(cpx_cpx_arbr7_fifo_rptr_a[1]), 
        .sel2(cpx_cpx_arbr7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel0), .psel1(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel1), .psel2(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel2), .psel3(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel3), .psel4(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel4), .psel5(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel5), .psel6(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel6), .psel7(
        cpx_cpx_arbr7_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl0_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl0_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl0_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl0_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl0_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl0_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl0_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl0_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl1_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl1_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl1_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl1_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl1_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl1_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl1_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl1_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl2_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl2_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl2_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl2_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl2_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl2_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl2_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl2_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl3_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl3_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl3_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl3_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl3_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl3_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl3_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl3_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl4_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl4_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl4_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl4_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl4_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl4_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl4_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl4_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl5_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl5_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl5_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl5_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl5_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl5_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl5_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl5_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl6_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl6_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl6_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl6_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl6_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl6_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl6_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl6_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl7_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl7_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl7_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl7_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl7_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl7_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl7_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl7_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl8_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbl8_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl8_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl8_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbl8_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbl8_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbl8_fifo_rptr_a[0]), .sel1(pcx_pcx_arbl8_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbl8_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbl8_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr0_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr0_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr0_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr0_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr0_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr0_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr0_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr0_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr0_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr1_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr1_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr1_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr1_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr1_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr1_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr1_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr1_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr1_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr2_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr2_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr2_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr2_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr2_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr2_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr2_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr2_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr2_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr3_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr3_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr3_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr3_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr3_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr3_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr3_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr3_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr3_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr4_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr4_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr4_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr4_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr4_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr4_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr4_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr4_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr4_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr5_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr5_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr5_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr5_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr5_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr5_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr5_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr5_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr5_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr6_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr6_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr6_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr6_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr6_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr6_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr6_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr6_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr6_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr7_ard_i_mux_fmem15_8_c0_0 ( .sel0(
        pcx_pcx_arbr7_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr7_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel0), .psel1(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel1), .psel2(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel2), .psel3(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel3), .psel4(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel4), .psel5(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel5), .psel6(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel6), .psel7(
        pcx_pcx_arbr7_ard_i_mux_fmem15_8_psel7) );
  cl_dp1_pdec8_8x pcx_pcx_arbr7_ard_i_mux_fmem7_0_c0_0 ( .sel0(
        pcx_pcx_arbr7_fifo_rptr_a[0]), .sel1(pcx_pcx_arbr7_fifo_rptr_a[1]), 
        .sel2(pcx_pcx_arbr7_fifo_rptr_a[2]), .test(1'b1), .psel0(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel0), .psel1(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel1), .psel2(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel2), .psel3(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel3), .psel4(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel4), .psel5(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel5), .psel6(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel6), .psel7(
        pcx_pcx_arbr7_ard_i_mux_fmem7_0_psel7) );
  cl_dp1_pdec4_8x pcx_pcx_arbr4_ard_i_mux_fifo_req_c0_0 ( .sel0(
        pcx_pcx_arbr4_fifo_read_select[0]), .sel1(
        pcx_pcx_arbr4_fifo_read_select[1]), .test(1'b1), .psel0(
        pcx_pcx_arbr4_ard_i_mux_fifo_req_psel0), .psel1(
        pcx_pcx_arbr4_ard_i_mux_fifo_req_psel1), .psel2(
        pcx_pcx_arbr4_ard_i_mux_fifo_req_psel2), .psel3(
        pcx_pcx_arbr4_ard_i_mux_fifo_req_psel3) );
  cl_dp1_pdec4_8x pcx_pcx_arbr5_ard_i_mux_fifo_req_c0_0 ( .sel0(
        pcx_pcx_arbr5_fifo_read_select[0]), .sel1(
        pcx_pcx_arbr5_fifo_read_select[1]), .test(1'b1), .psel0(
        pcx_pcx_arbr5_ard_i_mux_fifo_req_psel0), .psel1(
        pcx_pcx_arbr5_ard_i_mux_fifo_req_psel1), .psel2(
        pcx_pcx_arbr5_ard_i_mux_fifo_req_psel2), .psel3(
        pcx_pcx_arbr5_ard_i_mux_fifo_req_psel3) );
  cl_dp1_pdec4_8x pcx_pcx_arbr6_ard_i_mux_fifo_req_c0_0 ( .sel0(
        pcx_pcx_arbr6_fifo_read_select[0]), .sel1(
        pcx_pcx_arbr6_fifo_read_select[1]), .test(1'b1), .psel0(
        pcx_pcx_arbr6_ard_i_mux_fifo_req_psel0), .psel1(
        pcx_pcx_arbr6_ard_i_mux_fifo_req_psel1), .psel2(
        pcx_pcx_arbr6_ard_i_mux_fifo_req_psel2), .psel3(
        pcx_pcx_arbr6_ard_i_mux_fifo_req_psel3) );
  cl_dp1_pdec4_8x pcx_pcx_arbr7_ard_i_mux_fifo_req_c0_0 ( .sel0(
        pcx_pcx_arbr7_fifo_read_select[0]), .sel1(
        pcx_pcx_arbr7_fifo_read_select[1]), .test(1'b1), .psel0(
        pcx_pcx_arbr7_ard_i_mux_fifo_req_psel0), .psel1(
        pcx_pcx_arbr7_ard_i_mux_fifo_req_psel1), .psel2(
        pcx_pcx_arbr7_ard_i_mux_fifo_req_psel2), .psel3(
        pcx_pcx_arbr7_ard_i_mux_fifo_req_psel3) );
  cl_dp1_pdec4_8x pcx_pcx_arbr8_ard_i_mux_fifo_req_c0_0 ( .sel0(
        pcx_pcx_arbr8_fifo_read_select[0]), .sel1(
        pcx_pcx_arbr8_fifo_read_select[1]), .test(1'b1), .psel0(
        pcx_pcx_arbr8_ard_i_mux_fifo_req_psel0), .psel1(
        pcx_pcx_arbr8_ard_i_mux_fifo_req_psel1), .psel2(
        pcx_pcx_arbr8_ard_i_mux_fifo_req_psel2), .psel3(
        pcx_pcx_arbr8_ard_i_mux_fifo_req_psel3) );
  cl_dp1_muxbuff2_8x cpx_cpx_arbl0_ard_i_mux_reqmux_c0_0 ( .in0(n107079), 
        .in1(cpx_cpx_arbl0_fifo_req_sel_a), .out0(
        cpx_cpx_arbl0_ard_i_mux_reqmux_buffout0), .out1(
        cpx_cpx_arbl0_ard_i_mux_reqmux_buffout1) );
  cl_dp1_muxbuff2_8x pcx_pcx_arbr4_ard_i_mux_reqmux_c0_0 ( .in0(n107513), 
        .in1(pcx_pcx_arbr4_fifo_req_sel_a), .out0(
        pcx_pcx_arbr4_ard_i_mux_reqmux_buffout0), .out1(
        pcx_pcx_arbr4_ard_i_mux_reqmux_buffout1) );
  cl_dp1_muxbuff2_8x pcx_pcx_arbr5_ard_i_mux_reqmux_c0_0 ( .in0(n107521), 
        .in1(pcx_pcx_arbr5_fifo_req_sel_a), .out0(
        pcx_pcx_arbr5_ard_i_mux_reqmux_buffout0), .out1(
        pcx_pcx_arbr5_ard_i_mux_reqmux_buffout1) );
  cl_dp1_muxbuff2_8x pcx_pcx_arbr6_ard_i_mux_reqmux_c0_0 ( .in0(n107529), 
        .in1(pcx_pcx_arbr6_fifo_req_sel_a), .out0(
        pcx_pcx_arbr6_ard_i_mux_reqmux_buffout0), .out1(
        pcx_pcx_arbr6_ard_i_mux_reqmux_buffout1) );
  cl_dp1_muxbuff2_8x pcx_pcx_arbr7_ard_i_mux_reqmux_c0_0 ( .in0(n107537), 
        .in1(pcx_pcx_arbr7_fifo_req_sel_a), .out0(
        pcx_pcx_arbr7_ard_i_mux_reqmux_buffout0), .out1(
        pcx_pcx_arbr7_ard_i_mux_reqmux_buffout1) );
  cl_dp1_muxbuff2_8x pcx_pcx_arbr8_ard_i_mux_reqmux_c0_0 ( .in0(n107544), 
        .in1(pcx_pcx_arbr8_fifo_req_sel_a), .out0(
        pcx_pcx_arbr8_ard_i_mux_reqmux_buffout0), .out1(
        pcx_pcx_arbr8_ard_i_mux_reqmux_buffout1) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_fmem17_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_fmem17_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        cpx_cpx_arbl0_write_fifo_a[17]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_fmem16_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_fmem16_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        cpx_cpx_arbl0_write_fifo_a[16]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_fmem15_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_fmem15_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        cpx_cpx_arbl0_write_fifo_a[15]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_fmem14_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_fmem14_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        cpx_cpx_arbl0_write_fifo_a[14]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_fmem4_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_fmem4_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_arbr8_write_fifo_a[4]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_fmem3_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_fmem3_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_arbr8_write_fifo_a[3]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_fmem2_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_fmem2_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_arbr8_write_fifo_a[2]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_fmem1_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_fmem1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_arbr8_write_fifo_a[1]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_fmem0_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_fmem0_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(
        pcx_pcx_arbr8_write_fifo_a[0]), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_reqreg_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_reqreg_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_penc2_8x cpx_cpx_arbl0_ard_i_mux_atom_c0_0 ( .sel0(n171645), .psel0(
        cpx_cpx_arbl0_ard_i_mux_atom_psel0), .psel1(
        cpx_cpx_arbl0_ard_i_mux_atom_psel1) );
  cl_dp1_penc2_8x cpx_cpx_arbl1_ard_i_mux_atom_c0_0 ( .sel0(n171566), .psel0(
        cpx_cpx_arbl1_ard_i_mux_atom_psel0), .psel1(
        cpx_cpx_arbl1_ard_i_mux_atom_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr5_ard_i_mux_atom_c0_0 ( .sel0(n168039), .psel0(
        pcx_pcx_arbr5_ard_i_mux_atom_psel0), .psel1(
        pcx_pcx_arbr5_ard_i_mux_atom_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr6_ard_i_mux_atom_c0_0 ( .sel0(n167927), .psel0(
        pcx_pcx_arbr6_ard_i_mux_atom_psel0), .psel1(
        pcx_pcx_arbr6_ard_i_mux_atom_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr7_ard_i_mux_atom_c0_0 ( .sel0(n167815), .psel0(
        pcx_pcx_arbr7_ard_i_mux_atom_psel0), .psel1(
        pcx_pcx_arbr7_ard_i_mux_atom_psel1) );
  cl_dp1_penc2_8x pcx_pcx_arbr8_ard_i_mux_atom_c0_0 ( .sel0(n167703), .psel0(
        pcx_pcx_arbr8_ard_i_mux_atom_psel0), .psel1(
        pcx_pcx_arbr8_ard_i_mux_atom_psel1) );
  cl_dp1_l1hdr_8x cpx_cpx_arbl0_ard_i_dff_qual_atomic_d1_c0_0 ( .l1clk(
        cpx_cpx_arbl0_ard_i_dff_qual_atomic_d1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_l1hdr_8x pcx_pcx_arbr8_ard_i_dff_qual_atomic_d1_c0_0 ( .l1clk(
        pcx_pcx_arbr8_ard_i_dff_qual_atomic_d1_l1clk), .l2clk(l2clk), .se(
        pcx_pcx_dpa_pcx_dps8_tcu_scan_en_out_7_unused), .pce(1'b1), .pce_ov(
        pcx_pcx_dpa_pcx_dps8_tcu_pce_ov_out_7_unused), .stop(1'b0), .aclk(
        pcx_pcx_dpa_pcx_dps8_ccx_aclk_out_7_unused), .bclk(
        pcx_pcx_dpa_pcx_dps8_ccx_bclk_out_7_unused) );
  cl_dp1_rep_m6_32x trep0_i0_i11 ( .in(cpu_rep0_in[11]), .out(cpu_rep0_out[11]) );
  cl_dp1_rep_m6_32x trep0_i0_i10 ( .in(cpu_rep0_in[10]), .out(cpu_rep0_out[10]) );
  cl_dp1_rep_m6_32x trep0_i0_i9 ( .in(cpu_rep0_in[9]), .out(cpu_rep0_out[9])
         );
  cl_dp1_rep_m6_32x trep0_i0_i8 ( .in(cpu_rep0_in[8]), .out(cpu_rep0_out[8])
         );
  cl_dp1_rep_m6_32x trep0_i0_i7 ( .in(cpu_rep0_in[7]), .out(cpu_rep0_out[7])
         );
  cl_dp1_rep_m6_32x trep0_i0_i6 ( .in(cpu_rep0_in[6]), .out(cpu_rep0_out[6])
         );
  cl_dp1_rep_m6_32x trep0_i0_i5 ( .in(cpu_rep0_in[5]), .out(cpu_rep0_out[5])
         );
  cl_dp1_rep_m6_32x trep0_i0_i4 ( .in(cpu_rep0_in[4]), .out(cpu_rep0_out[4])
         );
  cl_dp1_rep_m6_32x trep0_i0_i3 ( .in(cpu_rep0_in[3]), .out(cpu_rep0_out[3])
         );
  cl_dp1_rep_m6_32x trep0_i0_i2 ( .in(cpu_rep0_in[2]), .out(cpu_rep0_out[2])
         );
  cl_dp1_rep_m6_32x trep0_i0_i1 ( .in(cpu_rep0_in[1]), .out(cpu_rep0_out[1])
         );
  cl_dp1_rep_m6_32x trep0_i0_i0 ( .in(cpu_rep0_in[0]), .out(cpu_rep0_out[0])
         );
  cl_dp1_rep_m6_32x trep0_i1_i11 ( .in(cpu_rep0_in[23]), .out(cpu_rep0_out[23]) );
endmodule

